-------------------------------------------------------------------------
-- Henry Duwe
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- mux2t1_N.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of an N-bit wide 2:1
-- mux using structural VHDL, generics, and generate statements.
--
--
-- NOTES:
-- 1/6/20 by H3::Created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity BarrelDecoder5_32 is
   generic(N : integer := 32); -- Generic of type integer for input/output data width. Default value is 32.
   port(
       i_WA         : in std_logic_vector(4 downto 0);
       o_OUT        : out std_logic_vector(N-1 downto 0));

end BarrelDecoder5_32;

architecture structural of BarrelDecoder5_32 is
begin 
   with i_WA select
   o_OUT <= "00000000000000000000000000000001" when "00001",
	    "00000000000000000000000000000011" when "00010",
	    "00000000000000000000000000000111" when "00011",
	    "00000000000000000000000000001111" when "00100",
	    "00000000000000000000000000011111" when "00101",
	    "00000000000000000000000000111111" when "00110",
	    "00000000000000000000000001111111" when "00111",
	    "00000000000000000000000011111111" when "01000",
	    "00000000000000000000000111111111" when "01001",
	    "00000000000000000000001111111111" when "01010",
	    "00000000000000000000011111111111" when "01011",
	    "00000000000000000000111111111111" when "01100",
	    "00000000000000000001111111111111" when "01101",
	    "00000000000000000011111111111111" when "01110",
	    "00000000000000000111111111111111" when "01111",
	    "00000000000000001111111111111111" when "10000",
	    "00000000000000011111111111111111" when "10001",
	    "00000000000000111111111111111111" when "10010",
	    "00000000000001111111111111111111" when "10011",
	    "00000000000011111111111111111111" when "10100",
	    "00000000000111111111111111111111" when "10101",
	    "00000000001111111111111111111111" when "10110",
	    "00000000011111111111111111111111" when "10111",
	    "00000000111111111111111111111111" when "11000",
	    "00000001111111111111111111111111" when "11001",
	    "00000011111111111111111111111111" when "11010",
	    "00000111111111111111111111111111" when "11011",
	    "00001111111111111111111111111111" when "11100",
	    "00011111111111111111111111111111" when "11101",
	    "00111111111111111111111111111111" when "11110",
	    "01111111111111111111111111111111" when "11111",
            "00000000000000000000000000000000" when others;
  
end structural;
